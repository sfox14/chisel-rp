// the dual-port LRAM Verilog below is adapted from Dan Strother's example:
// http://danstrother.com/2010/09/11/inferring-rams-in-fpgas/
// Removes a_wr: XST can not implement true dual port RAM in Distributed RAM

module DualPortLutRAM #(
    parameter DATA = 72,
    parameter ADDR = 10,
    parameter FNAME = "pe.mem"
) (
    input   wire               clk,
    // Port A
    input   wire                a_wr,
    input   wire    [ADDR-1:0]  a_addr,
    input   wire    [DATA-1:0]  a_din,
    output  reg     [DATA-1:0]  a_dout,
    // Port B
    input   wire                b_wr,
    input   wire    [ADDR-1:0]  b_addr,
    input   wire    [DATA-1:0]  b_din,
    output  reg     [DATA-1:0]  b_dout
);
// Shared memory
(* ram_style="distributed" *) reg [DATA-1:0] mem [(2**ADDR)-1:0];

initial
begin
    $readmemh(FNAME, mem);
end

// Port A
always @(posedge clk) begin
    a_dout      <= mem[a_addr];
    //if(a_wr) begin
    //    a_dout      <= a_din;
    //    mem[a_addr] <= a_din;
    //end
end
// Port B
always @(posedge clk) begin
    //b_dout      <= mem[b_addr];
    if(b_wr) begin
        b_dout      <= b_din;
        mem[b_addr] <= b_din;
    end
end
endmodule
